// module queue 
// import rv32i_types::*; #(
//     parameter       WIDTH = 32,
//     parameter       LENGTHEXP = 0
// )(
//     input   clk, rst,

//     input   logic   [WIDTH - 1: 0]  wdata,
//     input   logic   enqueue,

//     output  logic   [WIDTH - 1: 0]  rdata,
//     input  logic   dequeue,
    
//     output  logic   is_full,
//     output  logic   is_empty
// );